module Forwarding_Unit(
	input  alu_result, //value to forward which is available after ALU
	input  loadedData,  //value to forward which is available after RAM
	output forward0, //forward value to ALU input 0
	output forward1 //forward value to ALU input 1
);


endmodule