`timescale 1ns / 1ps
module test_singleCycleCPU;

SingleCycleCPU dut(
	.init(1)
);

endmodule